
// Copyright © 2024, Julian Scheffers, see LICENSE for more information

`timescale 1ns/1ps


